2
,110,130
,270,130
