5
Pin,50,200,500
Wire,260,530,300,530,0,2
Res,75,300,500
Wire,360,530,400,530,2,3
Ind,5,400,500
Wire,460,530,510,530,3,4
Cap,1,510,500
Wire,570,530,600,530,4,1
Pout,50,600,500
