3
Pin,50,200,500
Wire,260,530,300,530,0,1
Res,75,300,500
Wire,360,530,400,530,1,2
Pout,50,400,500

