8
Switch,50,100
Wire,110,120,140,120,0,4
Switch,50,120
Wire,110,140,140,140,1,4
Switch,50,160
Wire,110,180,140,180,2,6
Switch,50,180
Wire,110,200,140,200,3,6
AND,140,100
Wire,200,130,230,150,4,5
AND,230,130
Wire,290,160,330,160,5,7
OR,140,160
Wire,200,190,230,170,6,5
LED,330,140

